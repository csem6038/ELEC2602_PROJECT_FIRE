library verilog;
use verilog.vl_types.all;
entity Arithmetic_Logic_Unit_vlg_vec_tst is
end Arithmetic_Logic_Unit_vlg_vec_tst;
