library verilog;
use verilog.vl_types.all;
entity proc_vlg_vec_tst is
end proc_vlg_vec_tst;
