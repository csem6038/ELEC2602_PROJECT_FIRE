library verilog;
use verilog.vl_types.all;
entity controlunit_vlg_vec_tst is
end controlunit_vlg_vec_tst;
